package shared_pkg;
    int error_count;
    int correct_count;
    bit test_finished;
endpackage